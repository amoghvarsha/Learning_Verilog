module top_module 
( 
    input in, 
    output out 
);

    // The 'in' wire drive the 'out' wire continuously 
    assign out = in;

endmodule
